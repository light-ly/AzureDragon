package core;    

endpackage